// 337 TA Provided Lab 2 Testbench
// This code serves as a test bench for the 1 bit adder design 

`timescale 1ns / 100ps

module tb_adder_16bit
();
	// Define local parameters used by the test bench
	localparam NUM_INPUT_BITS			= 16;
	localparam NUM_OUTPUT_BITS		= NUM_INPUT_BITS + 1;
	localparam MAX_OUTPUT_BIT			= NUM_OUTPUT_BITS - 1;
	localparam NUM_TEST_BITS 			= (NUM_INPUT_BITS * 2) + 1;
	localparam MAX_TEST_BIT				= NUM_TEST_BITS - 1;
	localparam NUM_TEST_CASES 		= 100;
	localparam MAX_TEST_VALUE 		= NUM_TEST_CASES - 1;
	localparam TEST_A_BIT					= 0;
	localparam TEST_B_BIT					= NUM_INPUT_BITS;
	localparam TEST_CARRY_IN_BIT	= MAX_TEST_BIT;
	localparam TEST_SUM_BIT				= 0;
	localparam TEST_CARRY_OUT_BIT	= MAX_OUTPUT_BIT;
	localparam TEST_DELAY					= 10;
	
	// Declare Design Under Test (DUT) portmap signals
	
	reg	[NUM_INPUT_BITS-1:0] tb_a;
	reg	[NUM_INPUT_BITS-1:0] tb_b;
	reg	tb_carry_in;
	reg	[NUM_INPUT_BITS-1:0] tb_sum;
	reg	tb_carry_out;
        reg 	no_match = 0;
   
	
	// Declare test bench signals
	integer tb_case = 0;
	integer tb_test_case = 0;
	reg [MAX_TEST_BIT:0] tb_test_inputs;
	reg [MAX_OUTPUT_BIT:0] tb_expected_outputs;


        //reg [15:0] a;
        //reg [15:0] b;
  
   

   
	// DUT port map
       adder_16bit DUT(.a(tb_a), .b(tb_b), .carry_in(tb_carry_in), .sum(tb_sum), .overflow(tb_carry_out));
//	adder_16bit DUT(.a(a), .b(b), .carry_in(carry_in), .sum(sum), .overflow(carry_out));
	// Connect individual test input bits to a vector for easier testing
	//assign tb_a[NUM_INPUT_BITS-1:0]					= tb_test_inputs[15:0];
	//assign tb_b[NUM_INPUT_BITS-1:0]					= tb_test_inputs[31:16];
	//assign tb_carry_in	= tb_test_inputs[32];
	
	// Test bench process
	initial
	  begin
	      // Initialize test inputs for DUT
	/*	tb_test_inputs = 0;
		
		// Interative Exhaustive Testing Loop
		for(tb_test_case = 0; tb_test_case < NUM_TEST_CASES; tb_test_case = tb_test_case + 1)
		begin
			// Send test input to the design
			tb_test_inputs = tb_test_case[MAX_TEST_BIT:0];
			
			// Wait for a bit to allow this process to catch up with assign statements triggered
			// by test input assignment above
			#1;
			
			// Calculate the expected outputs
			tb_expected_outputs = tb_a + tb_b + tb_carry_in;
			
			// Wait for DUT to process the inputs
			#(TEST_DELAY - 1);
			
			// Check the DUT's Sum output value
			if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!", tb_test_case);
			end
			else
			begin
				$error("Incorrect Sum value for test case %d!", tb_test_case);
			end
			
			// Check the DUT's Carry Out output value
			if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!", tb_test_case);
			end
			else
			begin
				$error("Incorrect Carry Out value for test case %d!", tb_test_case);
			end
		end*/
	     //test case0
             tb_a = 16'b0000000000000000;
	     tb_b = 16'b0000000000000000;
	     no_match = 0;
	     
	     tb_carry_in = 1'b0;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			        no_match = 1;
			end
	     tb_case = tb_case + 1;
	     //test case1
             tb_a = 16'b1111111111111111;
	     tb_b = 16'b0000000000000001;
	     
	     tb_carry_in = 1'b0;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			   no_match = 1;
			   
			end
	     tb_case = tb_case + 1;
	     //test case2
	     tb_a = 16'b1111111111111111;
	     tb_b = 16'b1111111111111111;
	     no_match = 0;
	     
	     tb_carry_in = 1'b0;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			   no_match = 1;
			   
			end
	     tb_case = tb_case + 1;
              //test case1
	     tb_a = 16'b1010101010101010;
	     tb_b = 16'b0101010101010101;
	     no_match = 0;
	     
	     tb_carry_in = 1'b1;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			end
	     tb_case = tb_case + 1;
	   //test case 2
           tb_a = 16'b1010101010101010;
	     tb_b = 16'b0101010101010101;
	     no_match = 0;
	     
	     tb_carry_in = 1'b1;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			   no_match = 1;
			   
			end
	     tb_case = tb_case + 1;

            //test case 3
             tb_a = 16'b1111111111111111;
	     tb_b = 16'b0000000000000010;
	     no_match = 0;
	     
	     tb_carry_in = 1'b0;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			   no_match = 1;
			   
			end
	     tb_case = tb_case + 1;

	      //test case 4
             tb_a = 16'b0000000011111111;
	     tb_b = 16'b0000000011111111;
	     no_match = 0;
	     
	     tb_carry_in = 1'b1;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			   no_match = 1;
			   
			end
	     tb_case = tb_case + 1;
	      //test case 4
             tb_a = 16'b0000000011111111;
	     tb_b = 16'b0000000011111111;
	     no_match = 0;
	     
	     tb_carry_in = 1'b0;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Sum value for test case %d!",tb_case);
			end
			
			// Check the DUT's Carry Out output value
		if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!",tb_case);
			end
			else
			begin
				$info("Incorrect Carry Out value for test case %d!",tb_case);
			   no_match = 1;
			   
			end
	     tb_case = tb_case + 1;
/*
              //test case2
	     tb_a = 16'b1010101010101010;
	     tb_b = 16'b0101010101010101;
	     
	     tb_carry_in = 1'b1;
	     #1
	     tb_expected_outputs = tb_a + tb_b + tb_carry_in;
	     #9
	     if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!");
			end
			else
			begin
				$error("Incorrect Sum value for test case %d!");
			end
			
			// Check the DUT's Carry Out output value
			if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!");
			end
			else
			begin
				$error("Incorrect Carry Out value for test case %d!");
			end*/
end
/*	       
//*********************************************************************************	     
		// Initialize test inputs for DUT
		tb_test_inputs = 0;
		
		// Interative Exhaustive Testing Loop
		for(tb_test_case = 0; tb_test_case < NUM_TEST_CASES; tb_test_case = tb_test_case + 1)
		begin
			// Send test input to the design
			tb_test_inputs = tb_test_case[MAX_TEST_BIT:0];
			
			// Wait for a bit to allow this process to catch up with assign statements triggered
			// by test input assignment above
			#1;
			
			// Calculate the expected outputs
			tb_expected_outputs = tb_a + tb_b + tb_carry_in;
			
			// Wait for DUT to process the inputs
			#(TEST_DELAY - 1);
			
			// Check the DUT's Sum output value
			if(tb_expected_outputs[15:0] == tb_sum[15:0])
			begin
				$info("Correct Sum value for test case %d!", tb_test_case);
			end
			else
			begin
				$error("Incorrect Sum value for test case %d!", tb_test_case);
			end
			
			// Check the DUT's Carry Out output value
			if(tb_expected_outputs[16] == tb_carry_out)
			begin
				$info("Correct Carry Out value for test case %d!", tb_test_case);
			end
			else
			begin
				$error("Incorrect Carry Out value for test case %d!", tb_test_case);
			end
		end
	end
//8888888888888888888888888888888888888888888888888888888888888	
  */
	// Wrap-up process
/*	final
	begin
		if(NUM_TEST_CASES != tb_test_case)
		begin
			// Didn't run the test bench through all test cases
			$display("This test bench was not run long enough to execute all test cases. Please run this test bench for at least a total of %d ns", (NUM_TEST_CASES * TEST_DELAY));
		end
		else
		begin
			// Test bench was run to completion
			$display("This test bench has run to completion");
		end
	end*/
endmodule
