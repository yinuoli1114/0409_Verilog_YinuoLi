// $Id: $
// File name:   adder_16bit.sv
// Created:     9/11/2014
// Author:      Yinuo Li
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: 16-bit adder
module adder_16bit
(
	input wire [15:0] a,
	input wire [15:0] b,
	input wire carry_in,
	output wire [15:0] sum,
	output wire overflow
);

   always @ (a,b,carry_in)
    begin
      assert((a < 2**16)&&(a >= 0))
      else $error("Input a is incorrect");
      assert((b < 2**16)&&(b >= 0))
      else $error("Input a is incorrect");
      assert((carry_in == 1'b1)||(carry_in == 1'b0))
      else $error("Ipunt carry_in is not a digital logic value");
    end

adder_nbit #(16) IX (.a(a), .b(b), .carry_in(carry_in), .sum(sum), .overflow(overflow));

	// STUDENT: Fill in the correct port map with parameter override syntax for using your n-bit ripple carry adder design to be an 8-bit ripple carry adder design
endmodule
