library verilog;
use verilog.vl_types.all;
entity key_xor is
    port(
        data            : in     vl_logic_vector(47 downto 0);
        key             : in     vl_logic_vector(47 downto 0);
        \out\           : out    vl_logic_vector(47 downto 0)
    );
end key_xor;
