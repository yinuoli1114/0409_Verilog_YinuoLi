library verilog;
use verilog.vl_types.all;
entity tb_flex_stp_sr is
end tb_flex_stp_sr;
