library verilog;
use verilog.vl_types.all;
entity tb_scl_edge is
end tb_scl_edge;
