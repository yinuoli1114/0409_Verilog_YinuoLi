// $Id: $
// File name:   tb_key_xor.sv
// Created:     11/28/2014
// Author:      Jason Lin
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: testbench key xor
