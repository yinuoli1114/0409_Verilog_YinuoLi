// $Id: $
// File name:   tb_des_controller.sv
// Created:     11/19/2014
// Author:      Jason Lin
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Testbench for DES controller
