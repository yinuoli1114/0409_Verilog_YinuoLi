library verilog;
use verilog.vl_types.all;
entity des_2 is
    port(
        clk             : in     vl_logic;
        n_rst           : in     vl_logic;
        data_in         : in     vl_logic_vector(63 downto 0);
        key_in          : in     vl_logic_vector(63 downto 0);
        ready           : in     vl_logic;
        rw_mode         : in     vl_logic;
        data_out        : out    vl_logic_vector(63 downto 0);
        next_data       : out    vl_logic
    );
end des_2;
