library verilog;
use verilog.vl_types.all;
entity tb_moore is
end tb_moore;
