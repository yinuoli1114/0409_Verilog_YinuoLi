library verilog;
use verilog.vl_types.all;
entity tb_adder_16bit is
end tb_adder_16bit;
