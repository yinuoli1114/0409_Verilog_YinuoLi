library verilog;
use verilog.vl_types.all;
entity tb_flex_counter is
end tb_flex_counter;
