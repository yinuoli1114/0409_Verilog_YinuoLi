library verilog;
use verilog.vl_types.all;
entity main_controller is
    port(
        clk             : in     vl_logic;
        n_rst           : in     vl_logic;
        i2c_start       : in     vl_logic;
        i2c_stop        : in     vl_logic;
        i2c_rw          : in     vl_logic;
        data_ready      : in     vl_logic;
        next_data       : in     vl_logic;
        des_ready       : out    vl_logic;
        dir_io_sel      : out    vl_logic;
        ag_enable       : out    vl_logic;
        key_activate_key1: out    vl_logic;
        key_activate_key2: out    vl_logic
    );
end main_controller;
