// $Id: $
// File name:   i2c_slave.sv
// Created:     10/21/2014
// Author:      Yinuo Li
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: i2c_slave wrapper file

module i2c_slave
(
input wire clk,
 input wire n_rst,
 input wire scl,
 input wire sda_in,
 output wire sda_out,
 input wire write_enable,
 input wire [7:0] write_data,
 output wire fifo_empty,
 output wire fifo_full
 );
 wire rising_edge_found;
 wire falling_edge_found;
 wire [1:0] sda_mode;
 
 wire tx_out;
 wire tx_enable;
 //wire [7:0] tx_data;
 wire load_data;
 
 wire read_enable;
 wire [7:0] read_data;

 
 //wire [7:0] starting_byte;
 wire rw_mode;
 wire address_match;
 wire stop_found;
 wire start_found;
 
 wire rx_enable;
 wire [7:0] rx_data;
 
 wire byte_received;
 wire ack_prep;
 wire check_ack;
 wire ack_done;
  
 scl_edge SCL_EDGE
 (
 .clk(clk),
  .n_rst(n_rst),
  .scl(scl),
  .rising_edge_found(rising_edge_found),
  .falling_edge_found(falling_edge_found)
  );
  sda_sel SDA_SEL
  (
  .tx_out(tx_out),
   .sda_mode(sda_mode),
   .sda_out(sda_out)
   );
   tx_sr TX_SR
   (
   .clk(clk),
    .n_rst(n_rst),
    .tx_out(tx_out),
    .falling_edge_found(falling_edge_found),
    .tx_enable(tx_enable),
    .tx_data(read_data),
    .load_data(load_data)
    );
    tx_fifo TX_FIFO
    (
    .clk(clk),
     .n_rst(n_rst),
     .read_enable(read_enable),
     .write_enable(write_enable),
     .write_data(write_data),
     .read_data(read_data),
     .fifo_empty(fifo_empty),
     .fifo_full(fifo_full)
     );
     decode DECODE
     (
     .clk(clk),
      .n_rst(n_rst),
      .scl(scl),
      .sda_in(sda_in),
      .starting_byte(rx_data),
      .rw_mode(rw_mode),
      .address_match(address_match),
      .stop_found(stop_found),
      .start_found(start_found)
      );
      rx_sr RX_SR
      (
      .clk(clk),
       .n_rst(n_rst),
       .sda_in(sda_in),
       .rising_edge_found(rising_edge_found),
       .rx_enable(rx_enable),
       .rx_data(rx_data)
       );
       timer TIMER
       (
       .clk(clk),
	.n_rst(n_rst),
	.rising_edge_found(rising_edge_found),
	.falling_edge_found(falling_edge_found),
	.stop_found(stop_found),
	.start_found(start_found),
	.byte_received(byte_received),
	.ack_prep(ack_prep),
	.check_ack(check_ack),
	.ack_done(ack_done)
	);
	controller CONTROLLER
	(
	.clk(clk),
	 .n_rst(n_rst),
	 .stop_found(stop_found),
	 .start_found(start_found),
	 .byte_received(byte_received),
	 .ack_prep(ack_prep),
	 .check_ack(check_ack),
	 .ack_done(ack_done),
	 .rw_mode(rw_mode),
	 .address_match(address_match),
	 .sda_in(sda_in),
	 .rx_enable(rx_enable),
	 .tx_enable(tx_enable),
	 .read_enable(read_enable),
	 .sda_mode(sda_mode),
	 .load_data(load_data)
	 );
 endmodule
	 
      
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
