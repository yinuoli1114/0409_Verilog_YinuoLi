library verilog;
use verilog.vl_types.all;
entity tb_counter_wrapper is
end tb_counter_wrapper;
