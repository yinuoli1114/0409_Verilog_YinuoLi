// $Id: $
// File name:   key_permutation1.sv
// Created:     11/9/2014
// Author:      Yinuo Li
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: first permutation of the encryption key

module key_permutation1
  (
   input wire [63:0] k_o,
   output wire [55:0] kout
   );
   assign kout[0] = k_o[56];
   assign kout[1] = k_o[48];
   assign kout[2] = k_o[40];
   assign kout[3] = k_o[32];
   assign kout[4] = k_o[24];
   assign kout[5] = k_o[16];
   assign kout[6] = k_o[8];
   
   assign kout[7] = k_o[0];
   assign kout[8] = k_o[57];
   assign kout[9] = k_o[49];
   assign kout[10] = k_o[41];
   assign kout[11] = k_o[33];
   assign kout[12] = k_o[25];
   assign kout[13] = k_o[17];
   
   assign kout[14] = k_o[9];
   assign kout[15] = k_o[1];
   assign kout[16] = k_o[58];
   assign kout[17] = k_o[50];
   assign kout[18] = k_o[42];
   assign kout[19] = k_o[34];
   assign kout[20] = k_o[26];

   assign kout[21] = k_o[18];
   assign kout[22] = k_o[10];
   assign kout[23] = k_o[2];
   assign kout[24] = k_o[59];
   assign kout[25] = k_o[51];
   assign kout[26] = k_o[43];
   assign kout[27] = k_o[35];

   assign kout[28] = k_o[62];
   assign kout[29] = k_o[54];
   assign kout[30] = k_o[46];
   assign kout[31] = k_o[38];
   assign kout[32] = k_o[30];
   assign kout[33] = k_o[22];
   assign kout[34] = k_o[14];

   assign kout[35] = k_o[6];
   assign kout[36] = k_o[61];
   assign kout[37] = k_o[53];
   assign kout[38] = k_o[45];
   assign kout[39] = k_o[37];
   assign kout[40] = k_o[29];
   assign kout[41] = k_o[21];

   assign kout[42] = k_o[13];
   assign kout[43] = k_o[5];
   assign kout[44] = k_o[60];
   assign kout[45] = k_o[52];
   assign kout[46] = k_o[44];
   assign kout[47] = k_o[36];
   assign kout[48] = k_o[28];

   assign kout[49] = k_o[20];
   assign kout[50] = k_o[12];
   assign kout[51] = k_o[4];
   assign kout[52] = k_o[27];
   assign kout[53] = k_o[19];
   assign kout[54] = k_o[11];
   assign kout[55] = k_o[3];
 endmodule
 
   

   
   

   
