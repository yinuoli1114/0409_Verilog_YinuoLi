library verilog;
use verilog.vl_types.all;
entity tb_round_counter is
end tb_round_counter;
